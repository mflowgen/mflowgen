//-------------------------------------------------------------------------
// ProcXcel__ProcClass_ProcRTL__XcelClass_ChecksumXcelRTL.sv
//-------------------------------------------------------------------------
// This is the file that should be overwritten with PyMTL genenrated
// SystemVerilog of the processor and the null accelerator. You will need
// to copy ProcXcel__ProcClass_ProcRTL__XcelClass_NullXcelRTL.sv
// generated during Task 4.3 to overwrite this file. After making sure
// this file has the processor+accelerator to be pushed through the ASIC
// flow, you might also want to check that outputs/design.v indeed points
// to this file.
