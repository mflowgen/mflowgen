../pkgs/base/stdcells.lef