../pkgs/base/rtk-tech.lef