//------------------------------------------------------------------------
// ChecksumRTL.sv
//------------------------------------------------------------------------
// This is the file that should be overwritten with PyMTL genenrated
// SystemVerilog of the checksum unit. You will need to copy ChecksumRTL.sv
// generated during Task 2.6 to overwrite this file. After making sure
// this file has the checksum unit to be pushed through the ASIC flow, you
// might also want to check that outputs/design.v indeed points to this file.
